library verilog;
use verilog.vl_types.all;
entity ARQ_Lab1_vlg_vec_tst is
end ARQ_Lab1_vlg_vec_tst;
