library verilog;
use verilog.vl_types.all;
entity Registrador_4_bits_vlg_vec_tst is
end Registrador_4_bits_vlg_vec_tst;
