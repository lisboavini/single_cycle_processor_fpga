library verilog;
use verilog.vl_types.all;
entity Register_4_bits_vlg_vec_tst is
end Register_4_bits_vlg_vec_tst;
